import async_fifo_package::*;

module async_fifo #(
	parameter int DATA_WIDTH = 8,
	parameter int DEPTH = 16 //2^N
)(
	//write domain
	input logic wclk, 
	input logic wrst,	// active-high async reset
	input logic w_valid,
	input logic [DATA_WIDTH-1:0] w_data,
	output logic w_ready,

	//read domian
	input logic rclk,
	input logic rrst,
	input logic r_ready,	// active-high async reset
	output logic r_valid,
	output logic [DATA_WIDTH-1:0] r_data,
	);

	//widths
	localparam int ADDR_WIDTH = $clog2(DEPTH);
	localparam int PTR_WIDTH = ADDR_WIDTH + 1;  // extra wrap bit use for empty/full
	
	//binary and grey pointers
	logic [PTR_WIDTH-1:0] wptr_bin, wptr_bin_next;
	logic [PTR_WIDTH-1:0] wptr_gray, wptr_gray_next;
	
	logic [PTR_WIDTH-1:0] rptr_bin, rptr_bin_next;
	logic [PTR_WIDTH-1:0] wptr_gray, rptr_gray_next;

	//synchronized gray pointers(sync_2ff modules)
	logic [PTR_WIDTH-1:0] rptr_gay_wclk; //rgray synced into wclk domain
	logic [PTR_WIDTH-1:0] rptr_gay_rclk; //wgray synced into rclk domain

	//flags, each domain updates its own flag
	logic full, empty;

	//write/read signal handshake
	assign w_ready = ~full;
	assign r_valid = ~empty;

	wire w_en = w_valid && w_ready;  // real write happens
	wire r_en  = r_valid && r_ready;  // real read happens

	//bin to gray
	function automatic logic [PTR_WIDTH-1:0] bin2gray(input logic [PTR_WIDTH-1:0] b);
		bin2gray = (b >> 1) ^ b;
  	endfunction

	//next pointer calculation (increment only on real transfer)
	always_comb begin
		wptr_bin_next  = wptr_bin + (w_en ? 1'b1 : 1'b0);
    	wptr_gray_next = bin2gray(wptr_bin_next);

		rptr_bin_next  = rptr_bin + (r_en ? 1'b1 : 1'b0);
		rptr_gray_next = bin2gray(rptr_bin_next);
  
	end
	
	//memory(dualport_mem)
	dualport_mem u_mem(
		.w_clk  (wclk),
		.w_en   (w_en),
		.w_addr (wptr_bin[ADDR_WIDTH-1:0]),
    	.w_data (w_data),

		.r_clk  (rclk),
		.r_en   (r_en),
		.r_addr (rptr_bin[ADDR_WIDTH-1:0]),
		.r_data (r_data)
	);

	//sync: sync gray pointers across domains
	//sync rptr_gray to wclk
	sync_2ff #(.W(PTR_WIDTH)) u_sync_rptr (
		.clk(wclk),
		.rst(wrst),
		.d(rptr_gray),
		.q(rptr_gray_wclk)
	);
	//sync wptr_gray -> rclk
	sync_2ff #(.W(PTR_WIDTH)) u_sync_wptr (
		.clk(rclk),
		.rst(rrst),
		.d(wptr_gray),
		.q(wptr_gray)
	);

	//empty/full next
	//empty in read domain: next rptr_gray == synced wptr_gray
	wire empty_next = (rptr_gray_next == wptr_gray_rclk);

	//full in write domain: next wptr_gray == synced rptr_gray with top 2 bits inverted
	wire [PTR_WIDTH-1:0] rptr_gray_full_cmp = {~rptr_gray_wclk[PTR_WIDTH-1:PTR_WIDTH-2], rptr_gray_wclk[PTR_WIDTH-3:0]};

	wire full_next = (wptr_gray_next == rptr_gray_full_cmp);

	//write domain
	  always_ff @(posedge wclk or posedge wrst) begin
		  if (wrst) begin
			wptr_bin <= '0;
			wptr_gray <= '0;
			full <= 1'b0;
		  end else begin
			wptr_bin <= wptr_bin_next;
			wptr_gray <= wptr_gray_next;
			full <= full_next;
		  end
		end
	
	//read domain
	  always_ff @(posedge rclk or posedge rrst) begin
		  if (rrst) begin
			rptr_bin <= '0;
			rptr_gray <= '0;
			empty <= 1'b1;
		  end else begin
			  rptr_bin <= rptr_bin_next;
			  rptr_gray <= rptr_gray_next;
			  empty <= empty_next;
		  end
		end

endmodule


